----------------------------------------------------------------------
-- BCD mult 1x1 BCD
-- defines the memory content bit by bit.
-- C0 and D3 are simplified
----------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
Library UNISIM;
use UNISIM.vcomponents.all;

entity bcd_mul_mem2 is
    Port ( a : in  STD_LOGIC_VECTOR (3 downto 0);
           b : in  STD_LOGIC_VECTOR (3 downto 0);
           c : out  STD_LOGIC_VECTOR (3 downto 0);
           d : out  STD_LOGIC_VECTOR (3 downto 0));
end bcd_mul_mem2;

architecture Behavioral of bcd_mul_mem2 is
  type memFunc is array (0 to 255) of STD_LOGIC;
  constant fd2: std_logic_vector(0 to 255) := 
              "0000000000------0000000000------" & "0000000000------0000000000------" & 
              "0000000000------0000000011------" & "0000000111------0000001111------" & 
              "0000011111------0000011110------" & "--------------------------------" & 
              "--------------------------------" & "--------------------------------";
              
  constant fd1: std_logic_vector(0 to 255) := 
              "0000000000------0000000000------0000000000------0000000111------" & 
              "0000011111------0000111100------0000111000------0001110001------" & 
              "0001100011------0001100110--------------------------------------" & 
              "----------------------------------------------------------------";

  constant fd0: std_logic_vector(0 to 255) := 
              "0000000000------0000000000------0000011111------0000111000------" & 
              "0001100011------0011001100------0011011001------0010010010------" & 
              "0010100101------0010101010--------------------------------------" & 
              "----------------------------------------------------------------";

  constant fc3: std_logic_vector(0 to 255) := 
              "0000000000------0000000011------0000100001------0001001000------" & 
              "0010000100------0000000000------0001000010------0000100100------" & 
              "0100001000------0110000000--------------------------------------" & 
              "----------------------------------------------------------------";
              
  constant fc2: std_logic_vector(0 to 255) := 
              "0000000000------0000111100------0011000110------0010010011------" & 
              "0100101001------0101010101------0100101001------0110010010------" & 
              "0011000110------0001111000--------------------------------------" & 
              "----------------------------------------------------------------";

  constant fc1: std_logic_vector(0 to 255) := 
              "0000000000------0011001100------0101001010------0110100001------" & 
              "0001100011------0000000000------0110001100------0100001011------" & 
              "0010100101------0001100110--------------------------------------" & 
              "----------------------------------------------------------------";           
              
begin

  d(3) <= a(3) and b(3) and a(0) and b(0);
  d(2) <= fd2(conv_integer(a & b));
  d(1) <= fd1(conv_integer(a & b));
  d(0) <= fd0(conv_integer(a & b));

  c(3) <= fc3(conv_integer(a & b));
  c(2) <= fc2(conv_integer(a & b));
  c(1) <= fc1(conv_integer(a & b));
  c(0) <= a(0) and b(0);
  
end Behavioral;

