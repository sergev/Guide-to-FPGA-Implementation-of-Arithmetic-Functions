----------------------------------------------------------------------
-- BCD mult 1x1 BCD
-- defines the memory content as a 256x8 matrix
----------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
Library UNISIM;
use UNISIM.vcomponents.all;

entity bcd_mul_mem1 is
    Port ( a : in  STD_LOGIC_VECTOR (3 downto 0);
           b : in  STD_LOGIC_VECTOR (3 downto 0);
           c : out  STD_LOGIC_VECTOR (3 downto 0);
           d : out  STD_LOGIC_VECTOR (3 downto 0));
end bcd_mul_mem1;

architecture Behavioral of bcd_mul_mem1 is
  type memrom is array (0 to 255) of STD_LOGIC_VECTOR (7 downto 0);
  signal mrom: memrom := (
  "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", 
  "00000000", "00000000", "--------", "--------", "--------", "--------", "--------", "--------", 
  "00000000", "00000001", "00000010", "00000011", "00000100", "00000101", "00000110", "00000111", 
  "00001000", "00001001", "--------", "--------", "--------", "--------", "--------", "--------", 
  "00000000", "00000010", "00000100", "00000110", "00001000", "00010000", "00010010", "00010100", 
  "00010110", "00011000", "--------", "--------", "--------", "--------", "--------", "--------", 
  "00000000", "00000011", "00000110", "00001001", "00010010", "00010101", "00011000", "00100001", 
  "00100100", "00100111", "--------", "--------", "--------", "--------", "--------", "--------", 
  "00000000", "00000100", "00001000", "00010010", "00010110", "00100000", "00100100", "00101000", 
  "00110010", "00110110", "--------", "--------", "--------", "--------", "--------", "--------", 
  "00000000", "00000101", "00010000", "00010101", "00100000", "00100101", "00110000", "00110101", 
  "01000000", "01000101", "--------", "--------", "--------", "--------", "--------", "--------", 
  "00000000", "00000110", "00010010", "00011000", "00100100", "00110000", "00110110", "01000010", 
  "01001000", "01010100", "--------", "--------", "--------", "--------", "--------", "--------", 
  "00000000", "00000111", "00010100", "00100001", "00101000", "00110101", "01000010", "01001001", 
  "01010110", "01100011", "--------", "--------", "--------", "--------", "--------", "--------", 
  "00000000", "00001000", "00010110", "00100100", "00110010", "01000000", "01001000", "01010110", 
  "01100100", "01110010", "--------", "--------", "--------", "--------", "--------", "--------", 
  "00000000", "00001001", "00011000", "00100111", "00110110", "01000101", "01010100", "01100011", 
  "01110010", "10000001", "--------", "--------", "--------", "--------", "--------", "--------", 
  "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", --10
  "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
  "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", --11
  "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
  "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", --12
  "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
  "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", --13
  "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
  "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", --14
  "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------",
  "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------", --15
  "--------", "--------", "--------", "--------", "--------", "--------", "--------", "--------"
  );
  
  Signal cont: STD_LOGIC_VECTOR (7 downto 0);

begin
  
--  d <= mrom(conv_integer(a&b))(7 downto 4);
--  c <= mrom(conv_integer(a&b))(3 downto 0);
  cont <= mrom(conv_integer(a & b));
  d <= cont(7 downto 4);
  c <= cont(3 downto 0);
  
end Behavioral;

-----------------------------------------------------------------------------------------

